module mm_chain_dp(
    input

);
    
endmodule